
module switching_logic(
input wire [127:0][15:0] real_in,
input wire [127:0][15:0] complex_in,
input wire [3:0] state_select



);